*TL431 model from EDN magazine: March 15,1990, page 180-181
*Programmable Precision Reference pkg:TO-92 2,3,1. pkg:DIP8 6,1,8
*Connections
*             Anode
*             | Cathode
*             | | Reference
*             | | |
.SUBCKT TL431 2 3 1
*
*Reference input stage
Q1   3 1 10 QINPUT
RIN 10 2 500K
*
*Internal reference voltage
VR  20 2 DC 1.7791
RVR 20 2 1G
*
*Pole/Zero modeling
GM  0 30 10 20 1
RGM 30 0 1MEG
*Pole/Zeros: Pole 1= RGM & CP2, 10KHz
*            Pole 2= RP2 & CP2, 60KHz
*            Pole 3= CP1 & RZ1, 500KHz
*
CP1 30 40 15.9P
RZ1 40 0 20K
RP2 30 50 10MEG
CP2 50 0 0.265P
*Gain stage voltage clamp
DC  0 30 DCLAMP
*
*Output stage
GO  3 2 50 0 2.5U
DR  2 3 DNOM
*
.MODEL DNOM D(IS=100E-15 RS=7)
.MODEL DCLAMP D(IS=0.1)
.MODEL QINPUT NPN (BF=1 VAF=11.15)
.ENDS TL431



*OPTO FEDE
*NPN Optoisolator
*Connections
*                    LED Anode
*                    | LED Cathode
*                    | | Emitter
*                    | | | Collector
*                    | | | | Base
*                    | | | | |
.SUBCKT OPTOCOUPLER 1 2 4 5 6
C1 8 0 1nF
D1 9 2 LED
G1 5 6 8 0 1
VH1 1 9 0V
H1 7 0 VH1 1E-2
Q1 5 6 4 QNPN
R1 7 8 450
.MODEL LED D(IS=2.5E-12 RS=.75 CJO=3.5E-11 N=2)
.MODEL QNPN NPN(IS=3.33E-11 NF=1.35 CJC=4.74E-11 CJE=167E-12 TF=9.23E-10 TR=1.48E-7 BF=95 BR=10 IKF=.1 VAF=100)
.ENDS OPTOCOUPLER




******************************SIN USO************************************************
**************************************




* MODELO DEL LFX98
* AUTOR: FEDERICO [12-01-06]
* CONEXIONES:    POSITIVE POWER SUPPLY
*                | OS ADJ
*                | | IN
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | | HLD CAP
*                | | | | | | LREF
*                | | | | | | | L
*                | | | | | | | |
.SUBCKT LFX98    1 2 3 4 5 6 7 8
D1 9 11 DIODE
D2 11 9 DIODE
RF 11 5 30K
RH 6 10 300
SW 9 10 8 7 VSW OFF
XU1 10 5 1 4 5 TL08X
XU2 3 11 1 4 9 TL08X
.MODEL DIODE D(IS=2.55E-9 RS=0.042 N=1.75 TT=5.76E-6 CJO=1.85E-11 VJ=0.75 M=0.333 BV=100 IBV=1E-5)
.MODEL VSW SW(VT=1.4 VH=0 RON=1 ROFF=100E6)
.SUBCKT TL08X 1   2   3   4   5
C1   11 12 3.498E-12
C2    6  7 15E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
BGND 99  0 V=V(3)*.5 + V(4)*.5
BB    7 99 I=I(VB)*4.715E6 - I(VC)*5E6 + I(VE)*5E6 + I(VLP)*5E6 - I(VLN)*5E6
GA    6  0 11 12 282.8E-6
GCM   0  6 10 99 8.942E-9
ISS   3 10 DC 195E-6
HLIM 90  0 VLIM 1K
J1   11  2 10 JX
J2   12  1 10 JX
R2    6  9 100E3
RD1   4 11 3.536E3
RD2   4 12 3.536E3
RO1   8  5 150
RO2   7 99 150
RP    3  4 2.143E3
RSS  10 99 1.026E6
VB    9  0 DC 0
VC    3 53 DC 2.2
VE   54  4 DC 2.2
VLIM  7  8 DC 0
VLP  91  0 DC 25
VLN   0 92 DC 25
.MODEL DX D(IS=800E-18)
.MODEL JX PJF(IS=15E-12 BETA=270.1E-6 VTO=-1)
.ENDS TL08X
.ENDS LFX98




*Es el modelo de un transistor que le puedo cambiar el beta
.SUBCKT PNP C B E PARAMS: BETA=100
Q1 C B E QPNP
.MODEL QPNP PNP(BF={BETA})
.ENDS PNP

.SUBCKT NPN C B E PARAMS: BETA=100
Q2 C B E QNPN
.MODEL QNPN NPN(BF={BETA})
.ENDS NPN

.SUBCKT JFET-P D G S PARAMS: VT=2 BETA=2.5E-3
J3 D G S JP
.MODEL JP PJF(VTO={-VT} BETA={BETA})
.ENDS JFET-P

.SUBCKT JFET-N D G S PARAMS: VT=-2 BETA=2.5E-3
J4 D G S JN
.MODEL JN NJF(VTO={VT} BETA={BETA})
.ENDS JFET-N





.SUBCKT MPF102 D G S
J4 D G S JN

.MODEL JN NJF(
+ VTO=-3
+ BETA=1.304000e-03
+ LAMBDA=2.250000e-03
+ RD=1
+ RS=1
+ CGD=1.600000e-12
+ CGS=2.414000e-12
+ IS=33.570000e-15
+ KF=9.882000e-18)

*+ ISR=322.400000e-15
*+ ALPHA=311.7 VK=243.6
*+ M=.3622
*+ VTOTC=-2.500000e-03
*+ BETATCE=-0.5
.ENDS MPF102



