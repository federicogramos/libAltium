*Lo hice yo
*Transformador con 1 secundario
*Connections:
*                Vprim+
*                 | Vprim-
*                 | | Vsec+
*                 | | | Vsec-
*                 | | | |
.SUBCKT TRAFO1SEC 1 2 3 4 PARAMS: N2N1=1 RESPRIM=0.1 RESSEC=0.1 LPRIM=1u LSEC=1p LMAG=1m
E1 8 9 6 2 {N2N1}
VF1 4 9 0V
F1 6 2 VF1 {N2N1}
Lm 6 2 {LMAG}
LP 1 5 {LPRIM}
LS 7 3 {LSEC}
RP 5 6 {RESPRIM}
RS 8 7 {RESSEC}
.ENDS TRAFO1SEC

*Lo hice yo
*Transformador con 2 secundarios
*Connections:
*                 Pri+
*                 |   Pri-
*                 |   |   Sec1+
*                 |   |   |   Sec1-
*                 |   |   |   |   Sec2+
*                 |   |   |   |   |   Sec2-
*                 |   |   |   |   |   |
*                 |   |   |   |   |   |
*                 |   |   |   |   |   |
*                 |   |   |   |   |   |
.SUBCKT TRAFO2SEC 1   2   3   4   5   6  PARAMS: N2N1=1 N3N1=1 RPRI=0.1 RSEC=0.1 RTER=0.1 LPRI=1u LSEC=1u LTER=1u LMAG=5m
E1 10 11 7 2 {N2N1}
E2 13 14 7 2 {N3N1}
VF1 4 11 0V
F1 7 2 VF1 {N2N1}
VF2 6 14 0V
F2 7 2 VF2 {N3N1}
Lm 7 2 {LMAG}
LP 8 7 {LPRI}
LS 10 9 {LSEC}
LT 13 12 {LTER}
RP 1 8 {RPRI}
RS 9 3 {RSEC}
RT 12 5 {RTER}
.ENDS TRAFO2SEC











*********************************************************



