*************************************************************************************
*Agregado el 24-03-2010

.SUBCKT LM317/TI in adj out
* PEI 08/98 p62
J1 in out 4 JN
Q2 5 5 6 QPL .1
Q3 5 8 9 QNL .2
Q4 8 5 7 QPL .1
Q5 81 8 out QNL .2
Q6 out 81 10 QPL .2
Q7 12 81 13 QNL .2
*Q8 10 5 11 QPL .2
Q8 10A 5 11 QPL .2
Q9 14 12 10 QPL .2
Q10 16 5 17 QPL .2
Q11 16 14 15 QNL .2 OFF
Q12 out 20 16 QPL .2
Q13 in 19 20 QNL .2
Q14 19 5 18 QPL .2
Q15 out 21 19 QPL .2
Q16 21 22 16 QPL .2
Q17 21 out 24 QNL .2
Q18 22 22 16 QPL .2
Q19 22 out 241 QNL .2
Q20 out 25 16 QPL .2
Q21 25 26 out QNL .2
Q22A 35 35 in QPL .2
Q22B 16 35 in QPL .2
Q23 35 16 30 QNL .2
Q24A 27 40 29 QNL .2
Q24B 27 40 28 QNL .2
Q25 in 31 41 QNL 5
Q26 in 41 32 QNL 50
D1 out 4 DZ
D2 33 in DZ
D3 29 34 DZ
R1 in 6 310
R2 in 7 310
R3 in 11 190
R4 in 17 82
R5 in 18 5.6K
R6 4 8 100K
R7 8 81 130
*R8 10 12 12.4K
R8 10A 12 12.4K
R9 9 out 180
R10 13 out 4.1K
R11 14 out 5.8K
R12 15 out 72
R13 20 out 5.1K
R14 adj 24 12K
R15 24 241 2.4K
R16 16 25 6.7K
R17 16 40 12K
R18 30 41 130
R19 16 31 370
R20 26 27 13K
R21 27 40 400
R22 out 41 160
R23 33 34 18K
R24 28 29 160
R25 28 32 3
R26 32 out .1
C1 21 out 30PF
C2 21 adj 30PF
C3 25 26 5PF
CBS1 5 out 2PF
CBS2 35 out 1PF
CBS3 22 out 1PF
.MODEL JN NJF (BETA=1E-4 VTO=-7)
.MODEL DZ D(BV=6.3)
.MODEL QNL NPN (EG=1.22 BF=80 RB=100 CCS=1.5PF TF=.3NS TR=6NS
+ CJE=2PF CJC=1PF VAF=100 IS=1E-22 NF=1.2)
.MODEL QPL PNP (BF=40 RB=20 TF=.6NS TR=10NS CJE=1.5PF CJC=1PF VAF=50
+ IS=1E-22 NF=1.2)
.ENDS LM317/TI
*************************************************************************************




*Modelo UC3844
*Realizado por Federico Ramos
*24-02-08
*Pines para encapsulado DIP8
*              VFB  COMP    RT/CT  VREF GND VCC   ISENS OUTPUT
*              2    1       4      8    5   7     3     6
*              |    |       |      |    |   |     |     |
.SUBCKT UC3844 FEED EAOUTP  RTCT   REF  18  ALIM  VSEN  OUTP

*Node Bridge Data
ADVB1 [18 CLK REF REG SALCOMP][18$AD CLK$AD REF$AD REG$AD SALCOMP$AD] adc_mod
ADVB2 [REG$DA][REG] dac_mod
ADVB3 [6$DV NetFFT_4$DV QSAL$DV TOG$DV][6 NetFFT_4 QSAL TOG] dav_mod
.model adc_mod xadc
.model dac_mod xdac
.model dav_mod xdav

B2 ICOMPN 18 V=URAMP(V(11,18))-URAMP(V(11,18)-1)
B3 21 18 V=U(V(vsen,18)-V(icompn,18))*5
B6 ALIM 18 I=-I(BREF)
B8 5OA 18
+ V=U(V(TOG,18)-2.5)*U(V(REF,18)-2.5)*U(V(QSAL,18)-2.5)*U(V(CLK,18)-2.5)*10
BDISCH RTCT 18 I=(1-U(V(CLK,18)-2.5))*U(V(REG,18)-2.5)*(10/1000)
BREF REG 18 V=5*U(V(19,18)-6)
C1 18 6EA 15.9pF IC=0V
C2 18 3EA 200pF IC=0V
C5 18 2EA 0.02u IC=0V
CDELAY 18 SALCOMP 150pF IC=0V
CREF 18 REF 1nF IC=0V
D2 9 12 DIODO
D3 8OA 19 DIODO
D4 OUTP 8OA DIODO
D11 EAOUTP 12EA DIODO
D12 EAOUTP REF DIODO
D14 3EA 13EA DIODO
D15 18 6EA Di
E1 5EA 18 6EA 18 1
AFF [REG$AD 18$AD 18$AD SALCOMP$AD REF$AD CLK$AD][REG$DA QSAL$DV 6$DV]ffsrv2
AFFT [REG$AD 18$AD REF$AD CLK$AD][REG$DA TOG$DV NetFFT_4$DV]fft
G1 18 6EA 10EA FEED 100u
I2 REF EAOUTP 0.8mA
I3 19 8OA 100uA
I3EA 13EA 18 68uA
I4 18 1 0.9m
L1 2EA 3EA 10u
Q1 18 13EA 12EA PNPDEF
Q2 19 6OA OUTP NPNDEF
Q3 8OA 1 9OA NPNDEF
Q4 OUTP 9OA 18 NPNDEF
Q5 19 8OA 6OA NPNDEF
Q8 1 2OA 18 NPNDEF
R1 2OA 5OA 10K
R1EA 10EA REF 100K
R2 10EA 18 100K
R3 18 6EA 30meg
R4 12 11 2meg
R4EA 18 FEED 8meg
R6 11 18 1meg
R6EA 18 3EA 300
R7 VSEN 18 1meg
R9 2EA 5EA 5
RDELAY SALCOMP 21 1K
ROP REG 18 500
RPULL REF CLK 100K
RREG REG REF 0.33
RSTDBY ALIM 18 16.8K
RUVLO 19 18 1meg
SOSC CLK 18 RTCT 18 VSWOSC
SUVLO ALIM 19 ALIM 18 VSWUVLO
V4 EAOUTP 9 1V

.MODEL DIODO D()
.MODEL PNPDEF PNP()
.MODEL NPNDEF NPN()
.MODEL Di D(IS=1E-14 RS=1E+1 N=1E+0 TT=0E+0 CJO=0E+0 VJ=1E+0 M=5E-1 EG=1.11E+0 XTI=3E+0 KF=0E+0 AF=1E+0 FC=5E-1 BV=5E+0 IBV=1E-2)
.MODEL VSWOSC SW(VT=1.9E+0 VH=8.5E-1 RON=1E-2 ROFF=1E+6)
.MODEL VSWUVLO SW(VT=13 VH=3 RON=1E-2 ROFF=1E+6)
.MODEL ffsrv2 xsimcode(file="C:\FEDE\LIB_PROT\DIGITAL\ffsrv2.txt" func=ffsrv2)
.MODEL fft xsimcode(file="C:\FEDE\LIB_PROT\DIGITAL\fft.txt" func=fft)

.ENDS UC3844


*Del Protel (nombre original del modelo: AD620A)
* AD620A SPICE Macro-model              10/95, Rev. B
*                                       ARG / ADSC
*
* This version of the AD620 model simulates the worst-case
* parameters of the 'A' grade. The worst-case parameters
* used correspond to those in the data sheet.
*
*
* Revision History:
*     Rev. B
* Added V2,V3,V12,V13 and D3,D4,D15,D16 to clamp inputs to Q3,Q4 to
* prevent output phase reversal.
*
*
* Copyright 1990 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement. Use of this model
* indicates your acceptance with the terms and provisions in the License
* Statement.
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |  ref
*                |  |  |  |  |  |  rg1
*                |  |  |  |  |  |  |  rg2
*                |  |  |  |  |  |  |  |
.SUBCKT AD620    1  2  99 50 46 20 7  8
*
* INPUT STAGE
*
I1   7    50   5.002E-6
I2   8    50   5.002E-6
IOS  3    4    0.5E-9
VIOS 21   3    125E-6
CCM  3    4    2E-12
CD1  3    0    2E-12
CD2  4    0    2E-12
Q1   5    4    7    QN1
Q2   6    21   8    QN1
D1   7    4    DX
D2   8    21   DX
R1   1    3    400
R2   2    4    400
R3   99   5    100E3
R4   99   6    100E3
R5   7    9    24.7E3
R6   8    10   24.7E3
E1   9    46   11 5 375E6
E2   10   46   11 6 375E6
V1   99   11   0.5
RV1  99   11   1E3
CC1  5    9    4E-12
CC2  6    10   4E-12
*
* DIFFERENCE AMPLIFIER AND POLE AT 1MHZ
*
I3   18   50   5E-6
R7   99   12   11.937E3
R8   99   15   11.937E3
R9   14   18   1.592E3
R10  17   18   1.592E3
R11  9    13   10E3
R12  13   46   10E3
Q3   12   13   14   QN2
Q4   15   16   17   QN2
R13  19   16   10E3
R14  16   20   10E3
C1   12   15   6.667E-12
EOOS 19   10   POLY(1) (38,98) 1.5E-3 223.872
EREF 98   0    POLY(2) (99,0) (50,0) 0 0.5 0.5
D3 13 51 DX
D4 16 52 DX
V2 99 51 0.7
V3 99 52 0.7
D15 53 13 DX
D16 54 16 DX
V12 53 50 0.7
V13 54 50 0.7
*
* GAIN STAGE AND DOMINANT POLE AT 0.667HZ
*
R16  25   98   35.810E9
C2   25   98   6.667E-12
G1   98   25   12 15 83.776E-6
V6   99   26   1.53
V7   27   50   1.33
D7   25   26   DX
D8   27   25   DX
*
* POLE AT 10MHZ
*
R17  40   98   1
C3   40   98   15.916E-9
G2   98   40   25 98 1
*
* COMMON MODE STAGE WITH ZERO AT 708HZ
*
E3   36   98   POLY(2) (1,98) (2,98) 0 0.5 0.5
R18  36   38   1E6
R19  38   98   1
C5   36   38   224.812E-12
*
* OUTPUT STAGE
*
GSY  99   50   POLY(1) (99,50) 1.1725E-3 3.125E-6
RO1  99   45   250
RO2  45   50   250
L1   45   46   1E-6
GO1  45   99   99 40 4E-3
GO2  50   45   40 50 4E-3
GC1  43   50   40 45 4E-3
GC2  44   50   45 40 4E-3
F1   45   0    V4 1
F2   0    45   V5 1
V4   41   45   1.65
V5   45   42   1.65
D9   50   43   DY
D10  50   44   DY
D11  99   43   DX
D12  99   44   DX
D13  40   41   DX
D14  42   40   DX
*
* MODELS USED
*
.MODEL DX D(IS=1E-12)
.MODEL DY D(IS=1E-12 BV=50)
.MODEL QN1 NPN(BF=2.5E3 KF=0.7E-15 AF=1)
.MODEL QN2 NPN(BF=250 KF=0.5E-14 AF=1)
.ENDS AD620A

*************************************************************************************





